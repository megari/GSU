module gsu_mapper(
	input [23:0] addr,
	output [20:0] rom_addr,
	output is_rom,
	output [16:0] sram_addr,
	output is_sram
);



endmodule